library verilog;
use verilog.vl_types.all;
entity PRB_IB is
    port(
        Y               : out    vl_logic
    );
end PRB_IB;
