library verilog;
use verilog.vl_types.all;
entity DL2C_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end DL2C_UDP;
