`timescale 1 ns/100 ps
// Version: v11.5 SP2 11.5.2.6


module RAM_64_8_DP_RAM_64_8_DP_0_URAM(
       A_DOUT,
       B_DOUT,
       C_DIN,
       A_ADDR,
       B_ADDR,
       C_ADDR,
       A_CLK,
       B_CLK,
       C_CLK,
       C_WEN
    );
output [7:0] A_DOUT;
output [7:0] B_DOUT;
input  [7:0] C_DIN;
input  [5:0] A_ADDR;
input  [5:0] B_ADDR;
input  [5:0] C_ADDR;
input  A_CLK;
input  B_CLK;
input  C_CLK;
input  C_WEN;

    wire VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    RAM64x18 RAM_64_8_DP_RAM_64_8_DP_0_URAM_R0C0 (.A_DOUT({nc0, nc1, 
        nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, A_DOUT[7], A_DOUT[6], 
        A_DOUT[5], A_DOUT[4], A_DOUT[3], A_DOUT[2], A_DOUT[1], 
        A_DOUT[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, nc16, 
        nc17, nc18, nc19, B_DOUT[7], B_DOUT[6], B_DOUT[5], B_DOUT[4], 
        B_DOUT[3], B_DOUT[2], B_DOUT[1], B_DOUT[0]}), .BUSY(), 
        .A_ADDR_CLK(A_CLK), .A_DOUT_CLK(VCC), .A_ADDR_SRST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .A_ADDR_ARST_N(VCC), .A_DOUT_ARST_N(VCC), 
        .A_ADDR_EN(VCC), .A_DOUT_EN(VCC), .A_BLK({VCC, VCC}), .A_ADDR({
        GND, A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND, GND}), .B_ADDR_CLK(B_CLK), .B_DOUT_CLK(
        VCC), .B_ADDR_SRST_N(VCC), .B_DOUT_SRST_N(VCC), .B_ADDR_ARST_N(
        VCC), .B_DOUT_ARST_N(VCC), .B_ADDR_EN(VCC), .B_DOUT_EN(VCC), 
        .B_BLK({VCC, VCC}), .B_ADDR({GND, B_ADDR[5], B_ADDR[4], 
        B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND, GND}), 
        .C_CLK(C_CLK), .C_ADDR({GND, C_ADDR[5], C_ADDR[4], C_ADDR[3], 
        C_ADDR[2], C_ADDR[1], C_ADDR[0], GND, GND, GND}), .C_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, C_DIN[7], 
        C_DIN[6], C_DIN[5], C_DIN[4], C_DIN[3], C_DIN[2], C_DIN[1], 
        C_DIN[0]}), .C_WEN(C_WEN), .C_BLK({VCC, VCC}), .A_EN(VCC), 
        .A_ADDR_LAT(GND), .A_DOUT_LAT(VCC), .A_WIDTH({GND, VCC, VCC}), 
        .B_EN(VCC), .B_ADDR_LAT(GND), .B_DOUT_LAT(VCC), .B_WIDTH({GND, 
        VCC, VCC}), .C_EN(VCC), .C_WIDTH({GND, VCC, VCC}), .SII_LOCK(
        GND));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
