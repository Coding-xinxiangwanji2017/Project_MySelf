library verilog;
use verilog.vl_types.all;
entity CFG1_IP_B is
    port(
        IPB             : out    vl_logic;
        B               : in     vl_logic
    );
end CFG1_IP_B;
