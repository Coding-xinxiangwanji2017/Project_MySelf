library verilog;
use verilog.vl_types.all;
entity UDP_GBLAT is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end UDP_GBLAT;
