library verilog;
use verilog.vl_types.all;
entity PLL_V2 is
    generic(
        VCOFREQUENCY    : integer := 0;
        f_CLKA_LOCK     : integer := 3
    );
    port(
        CLKA            : in     vl_logic;
        EXTFB           : in     vl_logic;
        POWERDOWN       : in     vl_logic;
        OADIV0          : in     vl_logic;
        OADIV1          : in     vl_logic;
        OADIV2          : in     vl_logic;
        OADIV3          : in     vl_logic;
        OADIV4          : in     vl_logic;
        OAMUX0          : in     vl_logic;
        OAMUX1          : in     vl_logic;
        OAMUX2          : in     vl_logic;
        DLYGLA0         : in     vl_logic;
        DLYGLA1         : in     vl_logic;
        DLYGLA2         : in     vl_logic;
        DLYGLA3         : in     vl_logic;
        DLYGLA4         : in     vl_logic;
        OBDIV0          : in     vl_logic;
        OBDIV1          : in     vl_logic;
        OBDIV2          : in     vl_logic;
        OBDIV3          : in     vl_logic;
        OBDIV4          : in     vl_logic;
        OBMUX0          : in     vl_logic;
        OBMUX1          : in     vl_logic;
        OBMUX2          : in     vl_logic;
        DLYYB0          : in     vl_logic;
        DLYYB1          : in     vl_logic;
        DLYYB2          : in     vl_logic;
        DLYYB3          : in     vl_logic;
        DLYYB4          : in     vl_logic;
        DLYGLB0         : in     vl_logic;
        DLYGLB1         : in     vl_logic;
        DLYGLB2         : in     vl_logic;
        DLYGLB3         : in     vl_logic;
        DLYGLB4         : in     vl_logic;
        OCDIV0          : in     vl_logic;
        OCDIV1          : in     vl_logic;
        OCDIV2          : in     vl_logic;
        OCDIV3          : in     vl_logic;
        OCDIV4          : in     vl_logic;
        OCMUX0          : in     vl_logic;
        OCMUX1          : in     vl_logic;
        OCMUX2          : in     vl_logic;
        DLYYC0          : in     vl_logic;
        DLYYC1          : in     vl_logic;
        DLYYC2          : in     vl_logic;
        DLYYC3          : in     vl_logic;
        DLYYC4          : in     vl_logic;
        DLYGLC0         : in     vl_logic;
        DLYGLC1         : in     vl_logic;
        DLYGLC2         : in     vl_logic;
        DLYGLC3         : in     vl_logic;
        DLYGLC4         : in     vl_logic;
        FINDIV0         : in     vl_logic;
        FINDIV1         : in     vl_logic;
        FINDIV2         : in     vl_logic;
        FINDIV3         : in     vl_logic;
        FINDIV4         : in     vl_logic;
        FINDIV5         : in     vl_logic;
        FINDIV6         : in     vl_logic;
        FBDIV0          : in     vl_logic;
        FBDIV1          : in     vl_logic;
        FBDIV2          : in     vl_logic;
        FBDIV3          : in     vl_logic;
        FBDIV4          : in     vl_logic;
        FBDIV5          : in     vl_logic;
        FBDIV6          : in     vl_logic;
        FBDLY0          : in     vl_logic;
        FBDLY1          : in     vl_logic;
        FBDLY2          : in     vl_logic;
        FBDLY3          : in     vl_logic;
        FBDLY4          : in     vl_logic;
        FBSEL0          : in     vl_logic;
        FBSEL1          : in     vl_logic;
        XDLYSEL         : in     vl_logic;
        VCOSEL0         : in     vl_logic;
        VCOSEL1         : in     vl_logic;
        VCOSEL2         : in     vl_logic;
        GLA             : out    vl_logic;
        LOCK            : out    vl_logic;
        GLB             : out    vl_logic;
        YB              : out    vl_logic;
        GLC             : out    vl_logic;
        YC              : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of VCOFREQUENCY : constant is 1;
    attribute mti_svvh_generic_type of f_CLKA_LOCK : constant is 1;
end PLL_V2;
