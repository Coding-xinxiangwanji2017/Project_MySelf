library verilog;
use verilog.vl_types.all;
entity CMB7_primitive is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CMB7_primitive;
