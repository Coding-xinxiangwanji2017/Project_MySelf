library verilog;
use verilog.vl_types.all;
entity ABI_PLL_FRONT is
    generic(
        FB_MULTIPLIER   : integer := 1;
        VCOFREQUENCY    : real    := 0.000000
    );
    port(
        REFCK           : in     vl_logic;
        FB              : in     vl_logic;
        BYPASS          : in     vl_logic;
        RESET           : in     vl_logic;
        PD              : in     vl_logic;
        FSE             : in     vl_logic;
        MODE32K         : in     vl_logic;
        MODE_1V2        : in     vl_logic;
        MODE_3V3        : in     vl_logic;
        SSE             : in     vl_logic;
        DIVR5           : in     vl_logic;
        DIVR4           : in     vl_logic;
        DIVR3           : in     vl_logic;
        DIVR2           : in     vl_logic;
        DIVR1           : in     vl_logic;
        DIVR0           : in     vl_logic;
        RANGE3          : in     vl_logic;
        RANGE2          : in     vl_logic;
        RANGE1          : in     vl_logic;
        RANGE0          : in     vl_logic;
        DIVF9           : in     vl_logic;
        DIVF8           : in     vl_logic;
        DIVF7           : in     vl_logic;
        DIVF6           : in     vl_logic;
        DIVF5           : in     vl_logic;
        DIVF4           : in     vl_logic;
        DIVF3           : in     vl_logic;
        DIVF2           : in     vl_logic;
        DIVF1           : in     vl_logic;
        DIVF0           : in     vl_logic;
        DIVQ2           : in     vl_logic;
        DIVQ1           : in     vl_logic;
        DIVQ0           : in     vl_logic;
        SSMD1           : in     vl_logic;
        SSMD0           : in     vl_logic;
        SSMF4           : in     vl_logic;
        SSMF3           : in     vl_logic;
        SSMF2           : in     vl_logic;
        SSMF1           : in     vl_logic;
        SSMF0           : in     vl_logic;
        LOCKWIN2        : in     vl_logic;
        LOCKWIN1        : in     vl_logic;
        LOCKWIN0        : in     vl_logic;
        LOCKCNT3        : in     vl_logic;
        LOCKCNT2        : in     vl_logic;
        LOCKCNT1        : in     vl_logic;
        LOCKCNT0        : in     vl_logic;
        LOCK            : out    vl_logic;
        vco4x_normal    : out    vl_logic;
        vco4x_alt       : out    vl_logic;
        vco_000         : out    vl_logic;
        vco_000_alt     : out    vl_logic;
        vco_045         : out    vl_logic;
        vco_045_alt     : out    vl_logic;
        vco_090         : out    vl_logic;
        vco_090_alt     : out    vl_logic;
        vco_135         : out    vl_logic;
        vco_135_alt     : out    vl_logic;
        vco_180         : out    vl_logic;
        vco_180_alt     : out    vl_logic;
        vco_225         : out    vl_logic;
        vco_225_alt     : out    vl_logic;
        vco_270         : out    vl_logic;
        vco_270_alt     : out    vl_logic;
        vco_315         : out    vl_logic;
        vco_315_alt     : out    vl_logic;
        reset_reg       : out    vl_logic;
        divq_reset      : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of FB_MULTIPLIER : constant is 2;
    attribute mti_svvh_generic_type of VCOFREQUENCY : constant is 1;
end ABI_PLL_FRONT;
