library verilog;
use verilog.vl_types.all;
entity RCOSC is
    port(
        CLKOUT          : out    vl_logic
    );
end RCOSC;
