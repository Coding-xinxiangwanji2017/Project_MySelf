library verilog;
use verilog.vl_types.all;
entity CLKSRC is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end CLKSRC;
