library verilog;
use verilog.vl_types.all;
entity NVM is
    generic(
        MEMORYFILE      : string  := "";
        ACT_PROGFILE    : string  := "";
        ACT_CALIBRATIONDATA: integer := 0;
        FAST_SIM        : integer := 1;
        WR_THR          : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHK_CLK_RST     : integer := 0;
        RST_UNKNOWN     : integer := 1;
        POWERON_RESET   : integer := 2;
        CLK_UNKNOWN     : integer := 3;
        SAMPLE_CMD      : integer := 4;
        RD_DATA         : integer := 5;
        RD_LAST_WR      : integer := 6;
        COPY_PAGE_CA    : integer := 7;
        COPY_PAGE_CA1   : integer := 8;
        WR_DIFF_BLK     : integer := 9;
        WR_DIFF_BLK1    : integer := 10;
        WR_UPDATE_DATA  : integer := 11;
        WAIT_SP0_OVWR   : integer := 12;
        WAIT_SP0_OVWR1  : integer := 13;
        UPDATE_PG_CA    : integer := 14;
        UPDATE_PG_CA1   : integer := 15;
        PR_CHK_OVWRPRTC : integer := 16;
        RD_BLK_DLY      : integer := 17;
        RD_BLK_DLY1     : integer := 18;
        PR_OVWR_PROP    : integer := 19;
        PR_CHK_PROP     : integer := 20;
        RD_WAIT_CA      : integer := 21;
        RD_NEXT_BUSY    : integer := 22;
        DS_AB_INVALID   : integer := 23;
        ER_CHK_OVWRPRTC : integer := 24;
        ER_CHK_OVWRPRTC1: integer := 25;
        ER_AB_DLY       : integer := 26;
        ER_AB_DLY1      : integer := 27;
        UN_AB_PROP      : integer := 28;
        RD_WR_PIPE      : integer := 29;
        REMOVE_RESET    : integer := 30;
        RD_BLK_CA       : integer := 0;
        RD_BLK_CA1      : integer := 1;
        RD_DATA_CA      : integer := 2;
        RD_PIPE_DR      : integer := 3
    );
    port(
        ADDR            : in     vl_logic_vector(17 downto 0);
        WD              : in     vl_logic_vector(31 downto 0);
        DATAWIDTH       : in     vl_logic_vector(1 downto 0);
        REN             : in     vl_logic;
        READNEXT        : in     vl_logic;
        PAGESTATUS      : in     vl_logic;
        WEN             : in     vl_logic;
        ERASEPAGE       : in     vl_logic;
        PROGRAM         : in     vl_logic;
        SPAREPAGE       : in     vl_logic;
        AUXBLOCK        : in     vl_logic;
        UNPROTECTPAGE   : in     vl_logic;
        OVERWRITEPAGE   : in     vl_logic;
        DISCARDPAGE     : in     vl_logic;
        OVERWRITEPROTECT: in     vl_logic;
        PAGELOSSPROTECT : in     vl_logic;
        PIPE            : in     vl_logic;
        LOCKREQUEST     : in     vl_logic;
        CLK             : in     vl_logic;
        RESET           : in     vl_logic;
        RD              : out    vl_logic_vector(31 downto 0);
        BUSY            : out    vl_logic;
        STATUS          : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MEMORYFILE : constant is 1;
    attribute mti_svvh_generic_type of ACT_PROGFILE : constant is 1;
    attribute mti_svvh_generic_type of ACT_CALIBRATIONDATA : constant is 1;
    attribute mti_svvh_generic_type of FAST_SIM : constant is 1;
    attribute mti_svvh_generic_type of WR_THR : constant is 1;
    attribute mti_svvh_generic_type of CHK_CLK_RST : constant is 1;
    attribute mti_svvh_generic_type of RST_UNKNOWN : constant is 1;
    attribute mti_svvh_generic_type of POWERON_RESET : constant is 1;
    attribute mti_svvh_generic_type of CLK_UNKNOWN : constant is 1;
    attribute mti_svvh_generic_type of SAMPLE_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_DATA : constant is 1;
    attribute mti_svvh_generic_type of RD_LAST_WR : constant is 1;
    attribute mti_svvh_generic_type of COPY_PAGE_CA : constant is 1;
    attribute mti_svvh_generic_type of COPY_PAGE_CA1 : constant is 1;
    attribute mti_svvh_generic_type of WR_DIFF_BLK : constant is 1;
    attribute mti_svvh_generic_type of WR_DIFF_BLK1 : constant is 1;
    attribute mti_svvh_generic_type of WR_UPDATE_DATA : constant is 1;
    attribute mti_svvh_generic_type of WAIT_SP0_OVWR : constant is 1;
    attribute mti_svvh_generic_type of WAIT_SP0_OVWR1 : constant is 1;
    attribute mti_svvh_generic_type of UPDATE_PG_CA : constant is 1;
    attribute mti_svvh_generic_type of UPDATE_PG_CA1 : constant is 1;
    attribute mti_svvh_generic_type of PR_CHK_OVWRPRTC : constant is 1;
    attribute mti_svvh_generic_type of RD_BLK_DLY : constant is 1;
    attribute mti_svvh_generic_type of RD_BLK_DLY1 : constant is 1;
    attribute mti_svvh_generic_type of PR_OVWR_PROP : constant is 1;
    attribute mti_svvh_generic_type of PR_CHK_PROP : constant is 1;
    attribute mti_svvh_generic_type of RD_WAIT_CA : constant is 1;
    attribute mti_svvh_generic_type of RD_NEXT_BUSY : constant is 1;
    attribute mti_svvh_generic_type of DS_AB_INVALID : constant is 1;
    attribute mti_svvh_generic_type of ER_CHK_OVWRPRTC : constant is 1;
    attribute mti_svvh_generic_type of ER_CHK_OVWRPRTC1 : constant is 1;
    attribute mti_svvh_generic_type of ER_AB_DLY : constant is 1;
    attribute mti_svvh_generic_type of ER_AB_DLY1 : constant is 1;
    attribute mti_svvh_generic_type of UN_AB_PROP : constant is 1;
    attribute mti_svvh_generic_type of RD_WR_PIPE : constant is 1;
    attribute mti_svvh_generic_type of REMOVE_RESET : constant is 1;
    attribute mti_svvh_generic_type of RD_BLK_CA : constant is 1;
    attribute mti_svvh_generic_type of RD_BLK_CA1 : constant is 1;
    attribute mti_svvh_generic_type of RD_DATA_CA : constant is 1;
    attribute mti_svvh_generic_type of RD_PIPE_DR : constant is 1;
end NVM;
