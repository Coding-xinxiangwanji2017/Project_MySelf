library verilog;
use verilog.vl_types.all;
entity MACC_IP_P is
    port(
        clka            : in     vl_logic_vector(1 downto 0);
        a               : in     vl_logic_vector(17 downto 0);
        ea              : in     vl_logic_vector(1 downto 0);
        arsta_b         : in     vl_logic_vector(1 downto 0);
        srsta_b         : in     vl_logic_vector(1 downto 0);
        alat            : in     vl_logic_vector(1 downto 0);
        clkb            : in     vl_logic_vector(1 downto 0);
        b               : in     vl_logic_vector(17 downto 0);
        eb              : in     vl_logic_vector(1 downto 0);
        arstb_b         : in     vl_logic_vector(1 downto 0);
        srstb_b         : in     vl_logic_vector(1 downto 0);
        blat            : in     vl_logic_vector(1 downto 0);
        clkc            : in     vl_logic_vector(1 downto 0);
        c               : in     vl_logic_vector(43 downto 0);
        carryin         : in     vl_logic;
        ec              : in     vl_logic_vector(1 downto 0);
        arstc_b         : in     vl_logic_vector(1 downto 0);
        srstc_b         : in     vl_logic_vector(1 downto 0);
        clat            : in     vl_logic_vector(1 downto 0);
        cdin            : in     vl_logic_vector(43 downto 0);
        clksub          : in     vl_logic;
        sub             : in     vl_logic;
        esub            : in     vl_logic;
        alsub_b         : in     vl_logic;
        slsub_b         : in     vl_logic;
        sublat          : in     vl_logic;
        subad           : in     vl_logic;
        subsd_b         : in     vl_logic;
        clkshft         : in     vl_logic;
        shft            : in     vl_logic;
        eshft           : in     vl_logic;
        alshft_b        : in     vl_logic;
        slshft_b        : in     vl_logic;
        shftlat         : in     vl_logic;
        shftad          : in     vl_logic;
        shftsd_b        : in     vl_logic;
        clksel0         : in     vl_logic;
        sel0            : in     vl_logic;
        esel0           : in     vl_logic;
        alsel0_b        : in     vl_logic;
        slsel0_b        : in     vl_logic;
        sel0lat         : in     vl_logic;
        sel0ad          : in     vl_logic;
        sel0sd_b        : in     vl_logic;
        clksel1         : in     vl_logic;
        sel1            : in     vl_logic;
        esel1           : in     vl_logic;
        alsel1_b        : in     vl_logic;
        slsel1_b        : in     vl_logic;
        sel1lat         : in     vl_logic;
        sel1ad          : in     vl_logic;
        sel1sd_b        : in     vl_logic;
        clkp            : in     vl_logic_vector(1 downto 0);
        ep              : in     vl_logic_vector(1 downto 0);
        arstp_b         : in     vl_logic_vector(1 downto 0);
        srstp_b         : in     vl_logic_vector(1 downto 0);
        plat            : in     vl_logic_vector(1 downto 0);
        mode0           : in     vl_logic;
        mode1           : in     vl_logic;
        mode2           : in     vl_logic;
        pwrdwn_b        : in     vl_logic;
        p_out           : out    vl_logic_vector(43 downto 0);
        ovfl_ext_out    : out    vl_logic;
        cdout           : out    vl_logic_vector(43 downto 0)
    );
end MACC_IP_P;
