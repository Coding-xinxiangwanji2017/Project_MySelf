library verilog;
use verilog.vl_types.all;
entity CMEA_primitive is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CMEA_primitive;
