library verilog;
use verilog.vl_types.all;
entity ULSICC is
    port(
        LSICC           : in     vl_logic
    );
end ULSICC;
