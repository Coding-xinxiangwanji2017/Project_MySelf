library verilog;
use verilog.vl_types.all;
entity BUFF is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end BUFF;
