library verilog;
use verilog.vl_types.all;
entity FIFO4K18 is
    port(
        AEVAL11         : in     vl_logic;
        AEVAL10         : in     vl_logic;
        AEVAL9          : in     vl_logic;
        AEVAL8          : in     vl_logic;
        AEVAL7          : in     vl_logic;
        AEVAL6          : in     vl_logic;
        AEVAL5          : in     vl_logic;
        AEVAL4          : in     vl_logic;
        AEVAL3          : in     vl_logic;
        AEVAL2          : in     vl_logic;
        AEVAL1          : in     vl_logic;
        AEVAL0          : in     vl_logic;
        AFVAL11         : in     vl_logic;
        AFVAL10         : in     vl_logic;
        AFVAL9          : in     vl_logic;
        AFVAL8          : in     vl_logic;
        AFVAL7          : in     vl_logic;
        AFVAL6          : in     vl_logic;
        AFVAL5          : in     vl_logic;
        AFVAL4          : in     vl_logic;
        AFVAL3          : in     vl_logic;
        AFVAL2          : in     vl_logic;
        AFVAL1          : in     vl_logic;
        AFVAL0          : in     vl_logic;
        REN             : in     vl_logic;
        RBLK            : in     vl_logic;
        RCLK            : in     vl_logic;
        RESET           : in     vl_logic;
        RPIPE           : in     vl_logic;
        WEN             : in     vl_logic;
        WBLK            : in     vl_logic;
        WCLK            : in     vl_logic;
        RW2             : in     vl_logic;
        RW1             : in     vl_logic;
        RW0             : in     vl_logic;
        WW2             : in     vl_logic;
        WW1             : in     vl_logic;
        WW0             : in     vl_logic;
        ESTOP           : in     vl_logic;
        FSTOP           : in     vl_logic;
        WD17            : in     vl_logic;
        WD16            : in     vl_logic;
        WD15            : in     vl_logic;
        WD14            : in     vl_logic;
        WD13            : in     vl_logic;
        WD12            : in     vl_logic;
        WD11            : in     vl_logic;
        WD10            : in     vl_logic;
        WD9             : in     vl_logic;
        WD8             : in     vl_logic;
        WD7             : in     vl_logic;
        WD6             : in     vl_logic;
        WD5             : in     vl_logic;
        WD4             : in     vl_logic;
        WD3             : in     vl_logic;
        WD2             : in     vl_logic;
        WD1             : in     vl_logic;
        WD0             : in     vl_logic;
        RD17            : out    vl_logic;
        RD16            : out    vl_logic;
        RD15            : out    vl_logic;
        RD14            : out    vl_logic;
        RD13            : out    vl_logic;
        RD12            : out    vl_logic;
        RD11            : out    vl_logic;
        RD10            : out    vl_logic;
        RD9             : out    vl_logic;
        RD8             : out    vl_logic;
        RD7             : out    vl_logic;
        RD6             : out    vl_logic;
        RD5             : out    vl_logic;
        RD4             : out    vl_logic;
        RD3             : out    vl_logic;
        RD2             : out    vl_logic;
        RD1             : out    vl_logic;
        RD0             : out    vl_logic;
        FULL            : out    vl_logic;
        AFULL           : out    vl_logic;
        EMPTY           : out    vl_logic;
        AEMPTY          : out    vl_logic
    );
end FIFO4K18;
