library verilog;
use verilog.vl_types.all;
entity IO_DIFF is
    port(
        YIN             : in     vl_logic
    );
end IO_DIFF;
