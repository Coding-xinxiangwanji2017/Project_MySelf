library verilog;
use verilog.vl_types.all;
entity DLE2B_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end DLE2B_UDP;
