library verilog;
use verilog.vl_types.all;
entity INBUF_GTL25 is
    port(
        Y               : out    vl_logic;
        PAD             : in     vl_logic
    );
end INBUF_GTL25;
