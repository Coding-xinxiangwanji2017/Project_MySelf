library verilog;
use verilog.vl_types.all;
entity RCOSC_1MHZ is
    port(
        CLKOUT          : out    vl_logic
    );
end RCOSC_1MHZ;
