library verilog;
use verilog.vl_types.all;
entity MSSINT is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end MSSINT;
