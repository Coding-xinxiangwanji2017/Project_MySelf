library verilog;
use verilog.vl_types.all;
entity INBUF_HSTL_II is
    port(
        Y               : out    vl_logic;
        PAD             : in     vl_logic
    );
end INBUF_HSTL_II;
