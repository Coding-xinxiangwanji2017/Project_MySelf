library verilog;
use verilog.vl_types.all;
entity CCC_CONFIG is
    generic(
        CONFIG          : vl_logic_vector(209 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VCOFREQUENCY    : real    := 0.000000;
        WARNING_MSGS_ON : integer := 1
    );
    port(
        PCLK            : in     vl_logic;
        PRESET_N        : in     vl_logic;
        PSEL            : in     vl_logic;
        PWRITE          : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWDATA          : in     vl_logic_vector(7 downto 0);
        PADDR           : in     vl_logic_vector(7 downto 2);
        PRDATA          : out    vl_logic_vector(7 downto 0);
        CORE_LOCK       : in     vl_logic;
        RF_SEL          : out    vl_logic_vector(3 downto 0);
        RF_INV          : out    vl_logic;
        RF_DIV          : out    vl_logic_vector(7 downto 0);
        FB_SEL          : out    vl_logic_vector(3 downto 0);
        FB_INV          : out    vl_logic;
        FB_DIV          : out    vl_logic_vector(13 downto 0);
        GLMUX0_SEL      : out    vl_logic_vector(9 downto 0);
        GLMUX1_SEL      : out    vl_logic_vector(9 downto 0);
        GLMUX2_SEL      : out    vl_logic_vector(9 downto 0);
        GLMUX3_SEL      : out    vl_logic_vector(9 downto 0);
        GLMUX0_INV      : out    vl_logic;
        GLMUX1_INV      : out    vl_logic;
        GLMUX2_INV      : out    vl_logic;
        GLMUX3_INV      : out    vl_logic;
        GLMUX0_BUSY     : in     vl_logic;
        GLMUX1_BUSY     : in     vl_logic;
        GLMUX2_BUSY     : in     vl_logic;
        GLMUX3_BUSY     : in     vl_logic;
        GLMUX0_SELOUT   : out    vl_logic;
        GLMUX1_SELOUT   : out    vl_logic;
        GLMUX2_SELOUT   : out    vl_logic;
        GLMUX3_SELOUT   : out    vl_logic;
        GPD0_SEL        : out    vl_logic_vector(4 downto 0);
        GPD0_INV        : out    vl_logic;
        GPD0_DIV        : out    vl_logic_vector(7 downto 0);
        GPD0_NOPIPE_RSTSYNC: out    vl_logic;
        GPD1_SEL        : out    vl_logic_vector(4 downto 0);
        GPD1_INV        : out    vl_logic;
        GPD1_DIV        : out    vl_logic_vector(7 downto 0);
        GPD1_NOPIPE_RSTSYNC: out    vl_logic;
        GPD2_SEL        : out    vl_logic_vector(4 downto 0);
        GPD2_INV        : out    vl_logic;
        GPD2_DIV        : out    vl_logic_vector(7 downto 0);
        GPD2_NOPIPE_RSTSYNC: out    vl_logic;
        GPD3_SEL        : out    vl_logic_vector(4 downto 0);
        GPD3_INV        : out    vl_logic;
        GPD3_DIV        : out    vl_logic_vector(7 downto 0);
        GPD3_NOPIPE_RSTSYNC: out    vl_logic;
        GPD_SWRESYNC    : out    vl_logic;
        PLL_LOCKWIN     : out    vl_logic_vector(2 downto 0);
        PLL_LOCKCNT     : out    vl_logic_vector(3 downto 0);
        PLL_FBSEL       : out    vl_logic;
        PLL_SSE         : out    vl_logic;
        PLL_SSMD        : out    vl_logic_vector(1 downto 0);
        PLL_SSMF        : out    vl_logic_vector(4 downto 0);
        PLL_MODE_32K    : out    vl_logic;
        PLL_MODE_1V2    : out    vl_logic;
        PLL_MODE_3V3    : out    vl_logic;
        PLL_RANGE       : out    vl_logic_vector(3 downto 0);
        PLL_FBDIV       : out    vl_logic_vector(7 downto 0);
        PLL_CLKDIV      : out    vl_logic_vector(5 downto 0);
        PLL_VCODIV      : out    vl_logic_vector(2 downto 0);
        GPD0_G3STYLE_N  : out    vl_logic;
        GPD0_SRESETGENEN: out    vl_logic;
        GPD0_RESETGENEN : out    vl_logic;
        GPD1_G3STYLE_N  : out    vl_logic;
        GPD1_SRESETGENEN: out    vl_logic;
        GPD1_RESETGENEN : out    vl_logic;
        GPD2_G3STYLE_N  : out    vl_logic;
        GPD2_SRESETGENEN: out    vl_logic;
        GPD2_RESETGENEN : out    vl_logic;
        GPD3_G3STYLE_N  : out    vl_logic;
        GPD3_SRESETGENEN: out    vl_logic;
        GPD3_RESETGENEN : out    vl_logic;
        DELAY_LINE_SET  : out    vl_logic_vector(5 downto 0);
        DELAY_LINE_RF   : out    vl_logic;
        OVWR_SEL_RESET  : out    vl_logic;
        OVWR_VAL_RESET  : out    vl_logic;
        OVWR_SEL_PD     : out    vl_logic;
        OVWR_VAL_PD     : out    vl_logic;
        OVWR_SEL_BYPASS : out    vl_logic;
        OVWR_VAL_BYPASS : out    vl_logic;
        OVWR_SEL_GL     : out    vl_logic;
        OVWR_VAL_GL     : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CONFIG : constant is 2;
    attribute mti_svvh_generic_type of VCOFREQUENCY : constant is 1;
    attribute mti_svvh_generic_type of WARNING_MSGS_ON : constant is 1;
end CCC_CONFIG;
