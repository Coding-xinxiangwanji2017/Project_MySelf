library verilog;
use verilog.vl_types.all;
entity CLKINT is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end CLKINT;
