library verilog;
use verilog.vl_types.all;
entity CLKIO is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end CLKIO;
