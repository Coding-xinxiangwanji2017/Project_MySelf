library verilog;
use verilog.vl_types.all;
entity FCINIT_BUFF is
    port(
        FCO             : out    vl_logic;
        A               : in     vl_logic
    );
end FCINIT_BUFF;
