library verilog;
use verilog.vl_types.all;
entity CORERAM512X18 is
    generic(
        TC2CRWH         : integer := 503;
        TC2CWRH         : integer := 587;
        DYNAMIC         : integer := 1;
        MEMORYFILE      : string  := "";
        WARNING_MSGS_ON : integer := 1
    );
    port(
        RADDR8          : in     vl_logic;
        RADDR7          : in     vl_logic;
        RADDR6          : in     vl_logic;
        RADDR5          : in     vl_logic;
        RADDR4          : in     vl_logic;
        RADDR3          : in     vl_logic;
        RADDR2          : in     vl_logic;
        RADDR1          : in     vl_logic;
        RADDR0          : in     vl_logic;
        WADDR8          : in     vl_logic;
        WADDR7          : in     vl_logic;
        WADDR6          : in     vl_logic;
        WADDR5          : in     vl_logic;
        WADDR4          : in     vl_logic;
        WADDR3          : in     vl_logic;
        WADDR2          : in     vl_logic;
        WADDR1          : in     vl_logic;
        WADDR0          : in     vl_logic;
        RD17            : out    vl_logic;
        RD16            : out    vl_logic;
        RD15            : out    vl_logic;
        RD14            : out    vl_logic;
        RD13            : out    vl_logic;
        RD12            : out    vl_logic;
        RD11            : out    vl_logic;
        RD10            : out    vl_logic;
        RD9             : out    vl_logic;
        RD8             : out    vl_logic;
        RD7             : out    vl_logic;
        RD6             : out    vl_logic;
        RD5             : out    vl_logic;
        RD4             : out    vl_logic;
        RD3             : out    vl_logic;
        RD2             : out    vl_logic;
        RD1             : out    vl_logic;
        RD0             : out    vl_logic;
        WD17            : in     vl_logic;
        WD16            : in     vl_logic;
        WD15            : in     vl_logic;
        WD14            : in     vl_logic;
        WD13            : in     vl_logic;
        WD12            : in     vl_logic;
        WD11            : in     vl_logic;
        WD10            : in     vl_logic;
        WD9             : in     vl_logic;
        WD8             : in     vl_logic;
        WD7             : in     vl_logic;
        WD6             : in     vl_logic;
        WD5             : in     vl_logic;
        WD4             : in     vl_logic;
        WD3             : in     vl_logic;
        WD2             : in     vl_logic;
        WD1             : in     vl_logic;
        WD0             : in     vl_logic;
        RW1             : in     vl_logic;
        WW1             : in     vl_logic;
        RW0             : in     vl_logic;
        WW0             : in     vl_logic;
        REN             : in     vl_logic;
        RCLK            : in     vl_logic;
        WEN             : in     vl_logic;
        WCLK            : in     vl_logic;
        RESET           : in     vl_logic;
        PIPE            : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TC2CRWH : constant is 1;
    attribute mti_svvh_generic_type of TC2CWRH : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC : constant is 1;
    attribute mti_svvh_generic_type of MEMORYFILE : constant is 1;
    attribute mti_svvh_generic_type of WARNING_MSGS_ON : constant is 1;
end CORERAM512X18;
