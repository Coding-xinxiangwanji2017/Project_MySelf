library verilog;
use verilog.vl_types.all;
entity JKFFF is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end JKFFF;
