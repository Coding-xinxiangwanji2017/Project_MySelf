library verilog;
use verilog.vl_types.all;
entity IOINFF_BYPASS is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end IOINFF_BYPASS;
