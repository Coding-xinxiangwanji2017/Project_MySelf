library verilog;
use verilog.vl_types.all;
entity INV is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end INV;
