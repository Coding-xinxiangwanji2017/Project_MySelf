library verilog;
use verilog.vl_types.all;
entity CMEB_primitive is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CMEB_primitive;
