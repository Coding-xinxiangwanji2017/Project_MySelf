library verilog;
use verilog.vl_types.all;
entity DLN0 is
    port(
        G               : in     vl_logic;
        Q               : out    vl_logic;
        D               : in     vl_logic
    );
end DLN0;
