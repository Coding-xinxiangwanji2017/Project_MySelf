library verilog;
use verilog.vl_types.all;
entity DFN0 is
    port(
        CLK             : in     vl_logic;
        Q               : out    vl_logic;
        D               : in     vl_logic
    );
end DFN0;
