library verilog;
use verilog.vl_types.all;
entity DLN1C1 is
    port(
        CLR             : in     vl_logic;
        G               : in     vl_logic;
        Q               : out    vl_logic;
        D               : in     vl_logic
    );
end DLN1C1;
