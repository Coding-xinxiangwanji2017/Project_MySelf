library verilog;
use verilog.vl_types.all;
entity Dffpf is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end Dffpf;
