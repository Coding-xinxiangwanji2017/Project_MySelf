library verilog;
use verilog.vl_types.all;
entity CMA9_primitive is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CMA9_primitive;
