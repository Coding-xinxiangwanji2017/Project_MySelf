library verilog;
use verilog.vl_types.all;
entity IOIN_IB_ST is
    port(
        Y               : out    vl_logic;
        YIN             : in     vl_logic
    );
end IOIN_IB_ST;
