//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Apr 13 18:56:34 2016
// Version: v11.5 SP3 11.5.3.10
//////////////////////////////////////////////////////////////////////

`timescale 1 ns/100 ps

// RAM_2048_8_SDP
module RAM_2048_8_SDP(
    // Inputs
    RADDR,
    RCLK,
    REN,
    WADDR,
    WCLK,
    WD,
    WEN,
    // Outputs
    RD
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [10:0] RADDR;
input         RCLK;
input         REN;
input  [10:0] WADDR;
input         WCLK;
input  [7:0]  WD;
input         WEN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0]  RD;
//--------------------------------------------------------------------
// reg
//--------------------------------------------------------------------
reg [7:0]  RD_1;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [10:0] RADDR;
wire          RCLK;
wire   [7:0]  RD_0;
wire          REN;
wire   [10:0] WADDR;
wire          WCLK;
wire   [7:0]  WD;
wire          WEN;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire          GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign RD_0_net_0 = RD_0;
assign RD[7:0]    = RD_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------RAM_2048_8_SDP_RAM_2048_8_SDP_0_TPSRAM   -   Actel:SgCore:TPSRAM:1.0.101
RAM_2048_8_SDP_RAM_2048_8_SDP_0_TPSRAM RAM_2048_8_SDP_0(
        // Inputs
        .WD    ( WD ),
        .WADDR ( WADDR ),
        .RADDR ( RADDR ),
        .WEN   ( WEN ),
        .REN   ( REN ),
        .WCLK  ( WCLK ),
        .RCLK  ( RCLK ),
        // Outputs
        .RD    ( RD_0 ) 
        );
//register
always @(posedge RCLK)
begin
RD_1<=RD_0;
end

endmodule
