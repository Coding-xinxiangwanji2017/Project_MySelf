library verilog;
use verilog.vl_types.all;
entity IOOUTFF_BYPASS is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end IOOUTFF_BYPASS;
