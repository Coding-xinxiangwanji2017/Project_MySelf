library verilog;
use verilog.vl_types.all;
entity AB is
    generic(
        WIDTH           : integer := 32;
        MEMORYFILE      : string  := "";
        WARNING_MSGS_ON : integer := 1;
        ACT_DIE         : string  := "";
        ACT_PKG         : string  := "";
        FAST_ADC_CONV_SIM: integer := 0
    );
    port(
        VAREF           : inout  vl_logic;
        GNDREF          : in     vl_logic;
        AV0             : in     vl_logic;
        AC0             : in     vl_logic;
        AT0             : in     vl_logic;
        AV1             : in     vl_logic;
        AC1             : in     vl_logic;
        AT1             : in     vl_logic;
        AV2             : in     vl_logic;
        AC2             : in     vl_logic;
        AT2             : in     vl_logic;
        AV3             : in     vl_logic;
        AC3             : in     vl_logic;
        AT3             : in     vl_logic;
        AV4             : in     vl_logic;
        AC4             : in     vl_logic;
        AT4             : in     vl_logic;
        AV5             : in     vl_logic;
        AC5             : in     vl_logic;
        AT5             : in     vl_logic;
        AV6             : in     vl_logic;
        AC6             : in     vl_logic;
        AT6             : in     vl_logic;
        AV7             : in     vl_logic;
        AC7             : in     vl_logic;
        AT7             : in     vl_logic;
        AV8             : in     vl_logic;
        AC8             : in     vl_logic;
        AT8             : in     vl_logic;
        AV9             : in     vl_logic;
        AC9             : in     vl_logic;
        AT9             : in     vl_logic;
        ATRETURN01      : in     vl_logic;
        ATRETURN23      : in     vl_logic;
        ATRETURN45      : in     vl_logic;
        ATRETURN67      : in     vl_logic;
        ATRETURN89      : in     vl_logic;
        CMSTB0          : in     vl_logic;
        CMSTB1          : in     vl_logic;
        CMSTB2          : in     vl_logic;
        CMSTB3          : in     vl_logic;
        CMSTB4          : in     vl_logic;
        CMSTB5          : in     vl_logic;
        CMSTB6          : in     vl_logic;
        CMSTB7          : in     vl_logic;
        CMSTB8          : in     vl_logic;
        CMSTB9          : in     vl_logic;
        GDON0           : in     vl_logic;
        GDON1           : in     vl_logic;
        GDON2           : in     vl_logic;
        GDON3           : in     vl_logic;
        GDON4           : in     vl_logic;
        GDON5           : in     vl_logic;
        GDON6           : in     vl_logic;
        GDON7           : in     vl_logic;
        GDON8           : in     vl_logic;
        GDON9           : in     vl_logic;
        TMSTB0          : in     vl_logic;
        TMSTB1          : in     vl_logic;
        TMSTB2          : in     vl_logic;
        TMSTB3          : in     vl_logic;
        TMSTB4          : in     vl_logic;
        TMSTB5          : in     vl_logic;
        TMSTB6          : in     vl_logic;
        TMSTB7          : in     vl_logic;
        TMSTB8          : in     vl_logic;
        TMSTB9          : in     vl_logic;
        TMSTBINT        : in     vl_logic;
        DENAV0          : in     vl_logic;
        DENAC0          : in     vl_logic;
        DENAT0          : in     vl_logic;
        DENAV1          : in     vl_logic;
        DENAC1          : in     vl_logic;
        DENAT1          : in     vl_logic;
        DENAV2          : in     vl_logic;
        DENAC2          : in     vl_logic;
        DENAT2          : in     vl_logic;
        DENAV3          : in     vl_logic;
        DENAC3          : in     vl_logic;
        DENAT3          : in     vl_logic;
        DENAV4          : in     vl_logic;
        DENAC4          : in     vl_logic;
        DENAT4          : in     vl_logic;
        DENAV5          : in     vl_logic;
        DENAC5          : in     vl_logic;
        DENAT5          : in     vl_logic;
        DENAV6          : in     vl_logic;
        DENAC6          : in     vl_logic;
        DENAT6          : in     vl_logic;
        DENAV7          : in     vl_logic;
        DENAC7          : in     vl_logic;
        DENAT7          : in     vl_logic;
        DENAV8          : in     vl_logic;
        DENAC8          : in     vl_logic;
        DENAT8          : in     vl_logic;
        DENAV9          : in     vl_logic;
        DENAC9          : in     vl_logic;
        DENAT9          : in     vl_logic;
        MODE            : in     vl_logic_vector(3 downto 0);
        SYSCLK          : in     vl_logic;
        RTCCLK          : in     vl_logic;
        TVC             : in     vl_logic_vector(7 downto 0);
        STC             : in     vl_logic_vector(7 downto 0);
        VAREFSEL        : in     vl_logic;
        CHNUMBER        : in     vl_logic_vector(4 downto 0);
        ADCSTART        : in     vl_logic;
        PWRDWN          : in     vl_logic;
        ADCRESET        : in     vl_logic;
        ACMCLK          : in     vl_logic;
        ACMWEN          : in     vl_logic;
        ACMRESET        : in     vl_logic;
        ACMWDATA        : in     vl_logic_vector(7 downto 0);
        ACMADDR         : in     vl_logic_vector(7 downto 0);
        DAVOUT0         : out    vl_logic;
        DACOUT0         : out    vl_logic;
        DATOUT0         : out    vl_logic;
        DAVOUT1         : out    vl_logic;
        DACOUT1         : out    vl_logic;
        DATOUT1         : out    vl_logic;
        DAVOUT2         : out    vl_logic;
        DACOUT2         : out    vl_logic;
        DATOUT2         : out    vl_logic;
        DAVOUT3         : out    vl_logic;
        DACOUT3         : out    vl_logic;
        DATOUT3         : out    vl_logic;
        DAVOUT4         : out    vl_logic;
        DACOUT4         : out    vl_logic;
        DATOUT4         : out    vl_logic;
        DAVOUT5         : out    vl_logic;
        DACOUT5         : out    vl_logic;
        DATOUT5         : out    vl_logic;
        DAVOUT6         : out    vl_logic;
        DACOUT6         : out    vl_logic;
        DATOUT6         : out    vl_logic;
        DAVOUT7         : out    vl_logic;
        DACOUT7         : out    vl_logic;
        DATOUT7         : out    vl_logic;
        DAVOUT8         : out    vl_logic;
        DACOUT8         : out    vl_logic;
        DATOUT8         : out    vl_logic;
        DAVOUT9         : out    vl_logic;
        DACOUT9         : out    vl_logic;
        DATOUT9         : out    vl_logic;
        AG0             : out    vl_logic;
        AG1             : out    vl_logic;
        AG2             : out    vl_logic;
        AG3             : out    vl_logic;
        AG4             : out    vl_logic;
        AG5             : out    vl_logic;
        AG6             : out    vl_logic;
        AG7             : out    vl_logic;
        AG8             : out    vl_logic;
        AG9             : out    vl_logic;
        BUSY            : out    vl_logic;
        CALIBRATE       : out    vl_logic;
        DATAVALID       : out    vl_logic;
        SAMPLE          : out    vl_logic;
        RESULT          : out    vl_logic_vector(11 downto 0);
        RTCXTLMODE      : out    vl_logic_vector(1 downto 0);
        RTCXTLSEL       : out    vl_logic;
        RTCMATCH        : out    vl_logic;
        RTCPSMMATCH     : out    vl_logic;
        ACMRDATA        : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEMORYFILE : constant is 1;
    attribute mti_svvh_generic_type of WARNING_MSGS_ON : constant is 1;
    attribute mti_svvh_generic_type of ACT_DIE : constant is 1;
    attribute mti_svvh_generic_type of ACT_PKG : constant is 1;
    attribute mti_svvh_generic_type of FAST_ADC_CONV_SIM : constant is 1;
end AB;
