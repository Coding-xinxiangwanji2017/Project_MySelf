library verilog;
use verilog.vl_types.all;
entity IOENFF_BYPASS is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end IOENFF_BYPASS;
