library verilog;
use verilog.vl_types.all;
entity CMBB_primitive is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CMBB_primitive;
