library verilog;
use verilog.vl_types.all;
entity IO_UNUSED is
    port(
        YIN             : in     vl_logic;
        Y               : out    vl_logic
    );
end IO_UNUSED;
