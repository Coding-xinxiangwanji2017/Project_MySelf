library verilog;
use verilog.vl_types.all;
entity RCLKINT is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end RCLKINT;
